`include "src/simpleooo/param.v"

`include "src/simpleooo/cpu_ooo.v"

module top(
    input clk,
    input rst
);

reg init;
  always @(posedge clk) begin
    if (rst)
      init <= 1;
    else
      init <= 0;
   end


reg [`ROB_SIZE_LOG-1:0] ROB_tail_1, ROB_tail_2;
reg stall_1, stall_2, finish_1, finish_2, commit_deviation, addr_deviation, invalid_program;
reg C_mem_valid_r, C_mem_rdwt_r, C_is_br_r, C_taken_r;
reg [`MEMD_SIZE_LOG-1:0] C_mem_addr_r;


cpu_ooo copy1(.clk(stall_1 ? 0 : clk), .rst(rst));//, .C_valid(C_valid_1), .C_mem_valid(C_mem_valid_1), .C_mem_rdwt(C_mem_rdwt_1), .C_mem_addr(C_mem_addr_1), .C_is_br(C_is_br_1), .ROB_head(ROB_head_1), .ROB_tail(ROB_tail_1));
cpu_ooo copy2(.clk(stall_2 ? 0 : clk), .rst(rst));//, .C_valid(C_valid_2), .C_mem_valid(C_mem_valid_2), .C_mem_rdwt(C_mem_rdwt_2), .C_mem_addr(C_mem_addr_2), .C_is_br(C_is_br_2), .ROB_head(ROB_head_2), .ROB_tail(ROB_tail_2));

always @(posedge clk) begin
    if (rst) begin
        stall_1 <= 0;
        stall_2 <= 0;
        finish_1 <= 0;
        finish_2 <= 0;
        commit_deviation <= 0;
        invalid_program <= 0;
    end  
    else begin
    `ifndef IMM_STALL
        // If commit at same time, check if the program is valid
        if (!stall_1 && !stall_2 && copy1.C_valid && copy2.C_valid) begin
            if (copy1.C_mem_valid && copy1.C_mem_rdwt && copy2.C_mem_valid && copy2.C_mem_rdwt && (copy1.C_mem_addr == `SECRET_ADDR || copy2.C_mem_addr == `SECRET_ADDR))
                invalid_program <= 1;
        end
        else if (!stall_1 && !stall_2 && copy1.C_valid && !copy2.C_valid) begin
            stall_1 <= 1;
            commit_deviation <= 1;
            if (!(commit_deviation || ((`OBSV==`OBSV_EVERY_ADDR) ? addr_deviation : 0))) begin
                ROB_tail_1 <= copy1.ROB_tail;
                ROB_tail_2 <= copy2.ROB_tail;
            end
            // record the info of the early committed instruction
            C_mem_valid_r <= copy1.C_mem_valid;
            C_mem_rdwt_r <= copy1.C_mem_rdwt;
            C_mem_addr_r <= copy1.C_mem_addr;
            // C_is_br_r <= copy1.C_is_br;
            // C_taken_r <= copy1.C_taken;
        end
        else if (!stall_1 && !stall_2 && !copy1.C_valid && copy2.C_valid) begin
            stall_2 <= 1;
            commit_deviation <= 1;
            // Record the youngest instruction in ROB
            if (!commit_deviation) begin
                ROB_tail_1 <= copy1.ROB_tail;
                ROB_tail_2 <= copy2.ROB_tail;
            end
            C_mem_valid_r <= copy2.C_mem_valid;
            C_mem_rdwt_r <= copy2.C_mem_rdwt;
            C_mem_addr_r <= copy2.C_mem_addr;
            // C_is_br_r <= copy2.C_is_br;
            // C_taken_r <= copy2.C_taken;
        end
        // Compare the later committed instruction with the recorded early one
        else if (stall_1 && !stall_2 && copy2.C_valid) begin
            if (C_mem_valid_r && C_mem_rdwt_r && copy2.C_mem_valid && copy2.C_mem_rdwt && (C_mem_addr_r == `SECRET_ADDR || copy2.C_mem_addr == `SECRET_ADDR)) 
                invalid_program <= 1;
            // if (C_is_br_r && copy2.C_is_br && C_taken_r != copy2.C_taken)
            //     invalid_program <= 1;
            stall_1 <= 0;
        end
        else if (!stall_1 && stall_2 && copy1.C_valid) begin
            if (copy1.C_mem_valid && copy1.C_mem_rdwt && C_mem_valid_r && C_mem_rdwt_r && (C_mem_addr_r == `SECRET_ADDR || copy1.C_mem_addr == `SECRET_ADDR)) 
                invalid_program <= 1;
            // if (copy1.C_is_br && C_is_br_r && copy1.C_taken != C_taken_r)
            //     invalid_program <= 1;
            stall_2 <= 0;
        end
        `else
        if (!stall_1 && !stall_2 && copy1.C_valid && copy2.C_valid) begin
            if (copy1.C_mem_valid && copy1.C_mem_rdwt && copy2.C_mem_valid && copy2.C_mem_rdwt && ((`OBSV_LD_DATA) ? (copy1.C_rd_data!=copy2.C_rd_data): (copy1.C_mem_addr == `SECRET_ADDR || copy2.C_mem_addr == `SECRET_ADDR)))
                invalid_program = 1;
        end
        else if (!stall_1 && !stall_2 && copy1.C_valid && !copy2.C_valid) begin
            stall_1 = 1;
            commit_deviation <= 1;
            if (!(commit_deviation || ((`OBSV==`OBSV_EVERY_ADDR) ? addr_deviation : 0))) begin
                ROB_tail_1 <= copy1.ROB_tail;
                ROB_tail_2 <= copy2.ROB_tail;
            end
        end
        else if (!stall_1 && !stall_2 && !copy1.C_valid && copy2.C_valid) begin
            stall_2 = 1;
            commit_deviation <= 1;
            // Record the youngest instruction in ROB
            if (!(commit_deviation || ((`OBSV==`OBSV_EVERY_ADDR) ? addr_deviation : 0))) begin
                ROB_tail_1 <= copy1.ROB_tail;
                ROB_tail_2 <= copy2.ROB_tail;
            end
        end
        // Compare the later committed instruction with the recorded early one
        else if (stall_1 && !stall_2 && copy2.C_valid) begin
            if (copy1.C_mem_valid && copy1.C_mem_rdwt && copy2.C_mem_valid && copy2.C_mem_rdwt && ((`OBSV_LD_DATA) ? (copy1.C_rd_data!=copy2.C_rd_data): (copy1.C_mem_addr == `SECRET_ADDR || copy2.C_mem_addr == `SECRET_ADDR))) 
                invalid_program = 1;
            stall_1 <= 0;
        end
        else if (!stall_1 && stall_2 && copy1.C_valid) begin
            if (copy1.C_mem_valid && copy1.C_mem_rdwt && copy2.C_mem_valid && copy2.C_mem_rdwt && ((`OBSV_LD_DATA) ? (copy1.C_rd_data!=copy2.C_rd_data): (copy1.C_mem_addr == `SECRET_ADDR || copy2.C_mem_addr == `SECRET_ADDR))) 
                invalid_program = 1;
            stall_2 = 0;
        end
        `endif

        // Detect deviation in address (only consider this when no commit deviation has been found)
        if ((`OBSV==`OBSV_EVERY_ADDR) && !commit_deviation && copy1.ld_addr!=copy2.ld_addr) begin
            addr_deviation <= 1;
            ROB_tail_1 <= copy1.ROB_tail;
            ROB_tail_2 <= copy2.ROB_tail;
        end

        // Drain the ROB
        if ((commit_deviation || ((`OBSV==`OBSV_EVERY_ADDR) ? addr_deviation : 0)) && ((copy1.C_valid && copy1.ROB_head == ROB_tail_1-1 ) || (copy1.C_valid && copy1.C_squash)))
            finish_1 <= 1;
        if ((commit_deviation || ((`OBSV==`OBSV_EVERY_ADDR) ? addr_deviation : 0)) && ((copy2.C_valid && copy2.ROB_head == ROB_tail_1-1 ) || (copy2.C_valid && copy2.C_squash)))
            finish_2 <= 1;

        
    end
        

end



`ifdef INVARIANTS_FILE_1
    `include "scripts/induction_sandbox_2copy_SimpleOOO_DelayFuturistic/invariants.v"
`elsif INVARIANTS_FILE_2
    `include "scripts/induction_sandbox_2copy_SimpleOOO_noFwdFuturistic/invariants.v"
`else
    wire invariants = 1;
`endif

`define INDUCTION_K 20 // minimal 0, means no assumption at all
`define LOOK_AHEAD  20 // minimal 0, means no lookahead at all, i.e.,
                       // stop the simulation one cycle after K assumption finishes


// PART1: increment a counter
reg [10:0] counter;
always @(posedge clk) begin
    if (rst)
        counter <= 0;
    else if (counter <= (`INDUCTION_K + `LOOK_AHEAD))
        counter <= counter + 1;
end


// PART2: do assume in the first K cycle
reg [`LOOK_AHEAD:0] no_deviation_for_K;
always @(*)
    if (rst)
        no_deviation_for_K[0] = 1;
    else if (counter < `INDUCTION_K)
        if (commit_deviation || addr_deviation || !invariants)
            no_deviation_for_K[0] = 0;
        else
            no_deviation_for_K[0] = 1;
    else
        no_deviation_for_K[0] = 1;


// PART3: do assert in the K+1 cycle
reg [`LOOK_AHEAD:0] no_deviation_nextCycle;
always @(*)
    if (rst)
        no_deviation_nextCycle[0] = 1;
    else if (counter == `INDUCTION_K)
        if (commit_deviation || addr_deviation || !invariants)
            no_deviation_nextCycle[0] = 0;
        else
            no_deviation_nextCycle[0] = 1;
    else
        no_deviation_nextCycle[0] = 1;


// PART4: look ahead by simulating `LOOK_AHEAD more cycles
//        and check the assume and assert `LOOK_AHEAD cycles later
always @(posedge clk)
    if (`LOOK_AHEAD > 0)
        if (rst) begin
            no_deviation_for_K    [`LOOK_AHEAD:1] <= (1 << `LOOK_AHEAD) - 1;
            no_deviation_nextCycle[`LOOK_AHEAD:1] <= (1 << `LOOK_AHEAD) - 1;
        end else begin
            no_deviation_for_K    [`LOOK_AHEAD:1] <= no_deviation_for_K    [`LOOK_AHEAD-1:0];
            no_deviation_nextCycle[`LOOK_AHEAD:1] <= no_deviation_nextCycle[`LOOK_AHEAD-1:0];
        end

endmodule


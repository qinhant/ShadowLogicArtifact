// Step: Memory size. The instruction mem and data mem are stored in the same array
`define MEM_SIZE (`IMEM_SIZE + `DMEM_SIZE)
`define IMEM_SIZE 16
`define DMEM_SIZE 4

// Step: Regfile size and register length
`define RF_SIZE 4
`define REG_LEN 32